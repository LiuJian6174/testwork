1. main
2. jiliu
